`define SIZE 10
