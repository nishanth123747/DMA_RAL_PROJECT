`define SIZE 1
